module PWM_Generator_POWERTEST (
    input  i_clk, // 12MHz clock input 
    input  i_start, //button for start power test
    input  i_reset,
    output o_PWM_ESC, 
    output o_PWM_SERVO1, 
    output o_PWM_SERVO2
);

// module body 
//
    wire slow_clk_enable; // slow clock enable signal for debouncing FFs
    reg[27:0] counter_debounce=0;// counter for creating slow clock enable signals 
    wire tmp1,tmp2,duty_inc;// temporary flip-flop signals for debouncing the increasing button
    wire tmp3,tmp4,duty_dec;// temporary flip-flop signals for debouncing the decreasing button
//  counters for PWM output
    reg [18:0] counter_PWM_ESC; 
    reg [16:0] counter_PWM_SERVO1;
    reg [16:0] counter_PWM_SERVO2;


   //testing this change, will it set to 50% immediately?
   // reg[18:0] duty_cycle_Servo1 = 0;
   // reg[18:0] duty_cycle_Servo2 = 0;

   // normal values from working example
    reg[18:0] duty_cycle_Servo1 = 60000; 
    reg[16:0] duty_cycle_Servo2 = 60000; 
    reg[16:0] duty_cycle_ESC    = 6000; 


  // Debouncing 2 buttons for inc/dec duty cycle 
  // Firstly generate slow clock enable for debouncing flip-flop (4Hz)
 always @(posedge i_clk)
 begin
   counter_debounce <= counter_debounce + 1;
  
   //if(counter_debounce>=25000000) then  
   // for running on FPGA -- comment when running simulation

   if(counter_debounce>=1) 
   // for running simulation -- comment when running on FPGA
    counter_debounce <= 0;
 end
 // assign slow_clk_enable = counter_debounce == 25000000 ?1:0;
 // for running on FPGA -- comment when running simulation 

 assign slow_clk_enable = counter_debounce == 1 ? 1:0;


 // debouncing FFs for start  button  
 DFF_PWM PWM_DFF1(i_clk,slow_clk_enable,i_start,tmp1);
 DFF_PWM PWM_DFF2(i_clk,slow_clk_enable,tmp1, tmp2); 

 assign duty_inc =  tmp1 & (~ tmp2) & slow_clk_enable;



 // block  for on-off behavior
 always @(posedge i_clk) 
 begin
     if(i_reset == 0) begin
         duty_cycle_Servo1 <= 0; 
         duty_cycle_Servo2 <= 0;
         duty_cycle_ESC    <= 0;
     end
 // if button pressed
     else if (i_start == 1 && i_reset == 1) begin
         //set duty cycle to 50%
         //does the servo continuously move ? or do I have to send differing
         //signals? 
       //  duty_cycle_Servo1 <= duty_cycle_Servo1 + 12000; 
      //   duty_cycle_Servo2 <= duty_cycle_Servo1 + 12000;
       //  duty_cycle_ESC    <= duty_cycle_ESC    + 1200; 

	 duty_cycle_Servo1 <= 12000; 
         duty_cycle_Servo2 <= 12000;
         duty_cycle_ESC    <= 1200; 
     end   
 end         



 always @(posedge i_clk)
 begin 
   counter_PWM_SERVO1 <= counter_PWM_SERVO1 + 1; 
   if(counter_PWM_SERVO1 >= 240000)
       counter_PWM_SERVO1 <= 0; 
 end 
 assign o_PWM_SERVO1 = counter_PWM_SERVO1 < duty_cycle_Servo1 ? 1:0;
   
 always @(posedge i_clk)
 begin 
   counter_PWM_SERVO2 <= counter_PWM_SERVO2 + 1; 
   if(counter_PWM_SERVO2 >= 240000)
       counter_PWM_SERVO2 <= 0; 
 end 
 assign o_PWM_SERVO2 = counter_PWM_SERVO2 < duty_cycle_Servo2 ? 1:0;
 

 always @(posedge i_clk)
 begin
   counter_PWM_ESC <= counter_PWM_ESC + 1;
   if(counter_PWM_ESC>=24000) 
    counter_PWM_ESC <= 0;
 end
 assign o_PWM_ESC = counter_PWM_ESC < duty_cycle_ESC ? 1:0;
endmodule

module DFF_PWM(clk,en,D,Q);
input clk,en,D;
output reg Q;
always @(posedge clk)
begin 
 if(en==1) // slow clock enable signal 
  Q <= D;
end 
endmodule 

